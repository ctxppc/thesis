(
	do(
		pushScope
		set(abstract(cc.retcap), to: register(ra, cap(code)))
		set(abstract(ls.arg), to: 0)
		set(abstract(ls.arg$1), to: 1)
		set(register(a0), to: ls.arg)
		set(register(a1), to: ls.arg$1)
		call(capability(to: fib), parameters: a0 a1)
		set(abstract(df.result), to: register(a0, s32))
		set(register(a0), to: df.result)
		set(register(ra), to: cc.retcap)
		popScope
		return(to: register(ra, cap(code)))
	),
	procedures: (
		fib,
		in: do(
			pushScope
			set(abstract(cc.savedS1), to: register(s1, registerDatum))
			set(abstract(cc.savedS2), to: register(s2, registerDatum))
			set(abstract(cc.savedS3), to: register(s3, registerDatum))
			set(abstract(cc.savedS4), to: register(s4, registerDatum))
			set(abstract(cc.savedS5), to: register(s5, registerDatum))
			set(abstract(cc.savedS6), to: register(s6, registerDatum))
			set(abstract(cc.savedS7), to: register(s7, registerDatum))
			set(abstract(cc.savedS8), to: register(s8, registerDatum))
			set(abstract(cc.savedS9), to: register(s9, registerDatum))
			set(abstract(cc.savedS10), to: register(s10, registerDatum))
			set(abstract(cc.savedS11), to: register(s11, registerDatum))
			set(abstract(cc.retcap), to: register(ra, cap(code)))
			set(abstract(ls.first), to: register(a0, s32))
			set(abstract(ls.second), to: register(a1, s32))
			set(abstract(ls.arg), to: 2)
			set(abstract(ls.arg$1), to: 29)
			createVector(s32, count: 30, capability: abstract(ls.arg$2), scoped: false)
			set(register(a0), to: ls.arg)
			set(register(a1), to: ls.arg$1)
			set(register(a2), to: ls.arg$2)
			call(capability(to: recFib), parameters: a0 a1 a2)
			set(abstract(df.result$1), to: register(a0, s32))
			set(register(a0), to: df.result$1)
			set(register(s1), to: cc.savedS1)
			set(register(s2), to: cc.savedS2)
			set(register(s3), to: cc.savedS3)
			set(register(s4), to: cc.savedS4)
			set(register(s5), to: cc.savedS5)
			set(register(s6), to: cc.savedS6)
			set(register(s7), to: cc.savedS7)
			set(register(s8), to: cc.savedS8)
			set(register(s9), to: cc.savedS9)
			set(register(s10), to: cc.savedS10)
			set(register(s11), to: cc.savedS11)
			set(register(ra), to: cc.retcap)
			popScope
			return(to: register(ra, cap(code)))
		)
	)
	(
		recFib,
		in: do(
			pushScope
			set(abstract(cc.savedS1), to: register(s1, registerDatum))
			set(abstract(cc.savedS2), to: register(s2, registerDatum))
			set(abstract(cc.savedS3), to: register(s3, registerDatum))
			set(abstract(cc.savedS4), to: register(s4, registerDatum))
			set(abstract(cc.savedS5), to: register(s5, registerDatum))
			set(abstract(cc.savedS6), to: register(s6, registerDatum))
			set(abstract(cc.savedS7), to: register(s7, registerDatum))
			set(abstract(cc.savedS8), to: register(s8, registerDatum))
			set(abstract(cc.savedS9), to: register(s9, registerDatum))
			set(abstract(cc.savedS10), to: register(s10, registerDatum))
			set(abstract(cc.savedS11), to: register(s11, registerDatum))
			set(abstract(cc.retcap), to: register(ra, cap(code)))
			set(abstract(ls.index), to: register(a0, s32))
			set(abstract(ls.lastIndex), to: register(a1, s32))
			set(abstract(ls.nums), to: register(a2, cap(vector(of: s32, sealed: false))))
			if(
				do(
					set(abstract(ls.lhs), to: ls.index) set(abstract(ls.rhs), to: ls.lastIndex),
					then: relation(ls.lhs, gt, ls.rhs)
				),
				then: do(
					set(abstract(ls.vec), to: ls.nums)
					set(abstract(ls.idx), to: ls.lastIndex)
					getElement(of: abstract(ls.vec), index: ls.idx, to: abstract(df.result$2))
					set(register(a0), to: df.result$2)
					set(register(s1), to: cc.savedS1)
					set(register(s2), to: cc.savedS2)
					set(register(s3), to: cc.savedS3)
					set(register(s4), to: cc.savedS4)
					set(register(s5), to: cc.savedS5)
					set(register(s6), to: cc.savedS6)
					set(register(s7), to: cc.savedS7)
					set(register(s8), to: cc.savedS8)
					set(register(s9), to: cc.savedS9)
					set(register(s10), to: cc.savedS10)
					set(register(s11), to: cc.savedS11)
					set(register(ra), to: cc.retcap)
					popScope
					return(to: register(ra, cap(code)))
				),
				else: do(
					set(abstract(ls.vec$2), to: ls.nums)
					set(abstract(ls.idx$2), to: ls.index)
					set(abstract(ls.vec$3), to: ls.nums)
					set(abstract(ls.lhs$1), to: ls.index)
					set(abstract(ls.rhs$1), to: 2)
					compute(abstract(ls.idx$3), ls.lhs$1, sub, ls.rhs$1)
					getElement(of: abstract(ls.vec$3), index: ls.idx$3, to: abstract(ls.lhs$2))
					set(abstract(ls.vec$4), to: ls.nums)
					set(abstract(ls.lhs$3), to: ls.index)
					set(abstract(ls.rhs$2), to: 1)
					compute(abstract(ls.idx$4), ls.lhs$3, sub, ls.rhs$2)
					getElement(of: abstract(ls.vec$4), index: ls.idx$4, to: abstract(ls.rhs$3))
					compute(abstract(ls.elem$1), ls.lhs$2, add, ls.rhs$3)
					setElement(of: abstract(ls.vec$2), index: ls.idx$2, to: ls.elem$1)
					set(abstract(ls.lhs$4), to: ls.index)
					set(abstract(ls.rhs$4), to: 1)
					compute(abstract(ls.arg), ls.lhs$4, add, ls.rhs$4)
					set(abstract(ls.arg$1), to: ls.lastIndex)
					set(abstract(ls.arg$2), to: ls.nums)
					set(register(a0), to: ls.arg)
					set(register(a1), to: ls.arg$1)
					set(register(a2), to: ls.arg$2)
					call(capability(to: recFib), parameters: a0 a1 a2)
					set(abstract(df.result$3), to: register(a0, s32))
					set(register(a0), to: df.result$3)
					set(register(s1), to: cc.savedS1)
					set(register(s2), to: cc.savedS2)
					set(register(s3), to: cc.savedS3)
					set(register(s4), to: cc.savedS4)
					set(register(s5), to: cc.savedS5)
					set(register(s6), to: cc.savedS6)
					set(register(s7), to: cc.savedS7)
					set(register(s8), to: cc.savedS8)
					set(register(s9), to: cc.savedS9)
					set(register(s10), to: cc.savedS10)
					set(register(s11), to: cc.savedS11)
					set(register(ra), to: cc.retcap)
					popScope
					return(to: register(ra, cap(code)))
				)
			)
		)
	)
)