(
	do(
		pushScope()
		set(abstract(ls.arg0), to: constant(1))
		set(abstract(ls.arg1), to: constant(1))
		set(register(a0), to: abstract(ls.arg0))
		set(register(a1), to: abstract(ls.arg1))
		call(fib, parameters: a0 a1)
		set(abstract(df.result), to: register(a0, s32()))
		set(register(a0), to: abstract(df.result))
		popScope()
		return()
	),
	procedures: (
		fib,
		in: do(
			pushScope()
			set(abstract(ls.first), to: register(a0, s32()))
			set(abstract(ls.second), to: register(a1, s32()))
			set(abstract(ls.arg0), to: constant(2))
			set(abstract(ls.arg1), to: constant(29))
			pushVector(s32(), count: 30, into: abstract(ls.arg2))
			set(register(a0), to: abstract(ls.arg0))
			set(register(a1), to: abstract(ls.arg1))
			set(register(a2), to: abstract(ls.arg2))
			call(recFib, parameters: a0 a1 a2)
			set(abstract(df.result$1), to: register(a0, s32()))
			set(register(a0), to: abstract(df.result$1))
			popScope()
			return()
		)
	)
	(
		recFib,
		in: do(
			pushScope()
			set(abstract(ls.index), to: register(a0, s32()))
			set(abstract(ls.lastIndex), to: register(a1, s32()))
			set(abstract(ls.nums), to: register(a2, vectorCap(s32())))
			if(
				do(
					set(abstract(ls.lhs), to: abstract(ls.index)) set(abstract(ls.rhs), to: abstract(ls.lastIndex)),
					then: relation(abstract(ls.lhs), gt, abstract(ls.rhs))
				),
				then: do(
					set(abstract(ls.vec), to: abstract(ls.nums))
					set(abstract(ls.idx), to: abstract(ls.lastIndex))
					getElement(of: abstract(ls.vec), index: abstract(ls.idx), to: abstract(df.result$2))
					set(register(a0), to: abstract(df.result$2))
					popScope()
					return()
				),
				else: do(
					set(abstract(ls.lhs$1), to: abstract(ls.index))
					set(abstract(ls.rhs$1), to: constant(2))
					compute(abstract(ls.lhs$1), sub, abstract(ls.rhs$1), to: abstract(ls.indexOfFirst))
					set(abstract(ls.lhs$2), to: abstract(ls.index))
					set(abstract(ls.rhs$2), to: constant(1))
					compute(abstract(ls.lhs$2), sub, abstract(ls.rhs$2), to: abstract(ls.indexOfSecond))
					set(abstract(ls.lhs$3), to: abstract(ls.index))
					set(abstract(ls.rhs$3), to: constant(1))
					compute(abstract(ls.lhs$3), add, abstract(ls.rhs$3), to: abstract(ls.nextIndex))
					set(abstract(ls.vec$1), to: abstract(ls.nums))
					set(abstract(ls.idx$1), to: abstract(ls.indexOfFirst))
					getElement(of: abstract(ls.vec$1), index: abstract(ls.idx$1), to: abstract(ls.lhs$4))
					set(abstract(ls.vec$2), to: abstract(ls.nums))
					set(abstract(ls.idx$2), to: abstract(ls.indexOfSecond))
					getElement(of: abstract(ls.vec$2), index: abstract(ls.idx$2), to: abstract(ls.rhs$4))
					compute(abstract(ls.lhs$4), add, abstract(ls.rhs$4), to: abstract(ls.fibNum))
					set(abstract(ls.vec$3), to: abstract(ls.nums))
					set(abstract(ls.idx$3), to: abstract(ls.index))
					set(abstract(ls.elem), to: abstract(ls.fibNum))
					setElement(of: abstract(ls.vec$3), index: abstract(ls.idx$3), to: abstract(ls.elem))
					set(abstract(ls.arg0), to: abstract(ls.nextIndex))
					set(abstract(ls.arg1), to: abstract(ls.lastIndex))
					set(abstract(ls.arg2), to: abstract(ls.nums))
					set(register(a0), to: abstract(ls.arg0))
					set(register(a1), to: abstract(ls.arg1))
					set(register(a2), to: abstract(ls.arg2))
					call(recFib, parameters: a0 a1 a2)
					set(abstract(df.result$3), to: register(a0, s32()))
					set(register(a0), to: abstract(df.result$3))
					popScope()
					return()
				)
			)
		)
	)
)